`default_nettype none

`define     TRUE          1'b1
`define     FALSE         1'b0

`define     NULL          0
